module disp(

    );
endmodule
