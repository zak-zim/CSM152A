module tb();



endmodule
