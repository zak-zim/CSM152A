module StopTop();



endmodule
