module db();



endmodule