module StopController();



endmodule
