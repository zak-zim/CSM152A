module clock();


endmodule
