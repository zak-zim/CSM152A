module rps(move1, move2, result);

input move1;
input move2;
output result;

parameter ROCK = 2'b00;
parameter PAPER = 2'b01;
parameter SCISSORS = 2'b10;

endmodule