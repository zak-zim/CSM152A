module clock(

    );
endmodule
