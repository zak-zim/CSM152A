module StopTop(reset, clk, sel, adj, pause);

input reset;
input clk;
input sel;
input adj;
input pause;

reg counterClk;
reg adjClk;
reg dispClk;
reg blinkClk;
wire [2:0] enables;
wire [5:0] min;
wire [5:0] sec;

clock clock(clk, counterClk, adjClk, dispClk, blinkClk);
StopController controller(clk, adj, pause, enables);

endmodule
