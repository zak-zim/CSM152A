module ExtractLeadingBits(
input [11:0] dec, output [3:4] mant, output xBit
);

endmodule